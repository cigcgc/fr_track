`define MODULE_NAME FP_Sqrt_Top
`define NO_CE
