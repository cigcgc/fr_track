parameter DIN_WIDTH = 12;
parameter COEFF_WIDTH = 16;
parameter DOUT_WIDTH = 27;
parameter NUM_CHN = 1;
parameter NUM_FACTOR = 2;
parameter TAPS_SIZE = 128;
parameter NUM_TDM = 1;
parameter COEFF_PATH = "./coeff.dat";
