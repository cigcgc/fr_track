`define module_name CORDIC_Top2
`define VECTOR
`define PIPELINE
`define DEGREE_8_8
`define XY_BITS 17
`define THETA_BITS 17
`define ITERATIONS 16
`define ITERATION_BITS 4
