//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2A-LV18EQ144C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Tue Jun 20 11:13:56 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [10:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [28:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h64615E5B5855524F4B4845423F3C3935322F2C2926231F1C191613100D090603;
defparam prom_inst_0.INIT_RAM_01 = 256'hC8C5C2BFBCB8B5B2AFACA9A6A3A09D999693908D8A8784817D7A7774716E6B68;
defparam prom_inst_0.INIT_RAM_02 = 256'h292623201D1A1714110E0B080502FFFCF9F6F3F0EDEAE7E4E0DDDAD7D4D1CECB;
defparam prom_inst_0.INIT_RAM_03 = 256'h8885827F7C797774716E6B6865625F5C595653504D4A4744413E3B3835322F2C;
defparam prom_inst_0.INIT_RAM_04 = 256'hE3E0DDDBD8D5D2CFCDCAC7C4C1BFBCB9B6B3B0ADABA8A5A29F9C999794918E8B;
defparam prom_inst_0.INIT_RAM_05 = 256'h393734312F2C292724211F1C191714110F0C09070401FEFCF9F6F3F1EEEBE8E6;
defparam prom_inst_0.INIT_RAM_06 = 256'h74737271706F6E6D6C6B6A696867666562605D5B585653504E4B494644413E3C;
defparam prom_inst_0.INIT_RAM_07 = 256'hD4D2D0CECBC9C7C5C2C0BEBCB9B7B5B2B0AEABA9A7A4A29F908A857F7A787675;
defparam prom_inst_0.INIT_RAM_08 = 256'h18161412100E0C0A08060401FFFDFBF9F7F5F3F1EFECEAE8E6E4E2DFDDDBD9D7;
defparam prom_inst_0.INIT_RAM_09 = 256'h5452504E4D4B4947454442403E3C3A39373533312F2D2B2928262422201E1C1A;
defparam prom_inst_0.INIT_RAM_0A = 256'h8786848381807E7D7B7A7877757372706F6D6B6A6866656361605E5C5B595755;
defparam prom_inst_0.INIT_RAM_0B = 256'hB2B1B0AFADACABAAA8A7A6A5A3A2A19F9E9D9B9A989796949391908F8D8C8A89;
defparam prom_inst_0.INIT_RAM_0C = 256'hD3D2D1D0CFCECDCCCBCAC9C8C7C6C5C4C3C2C1C0BFBEBDBCBBBAB9B8B7B6B5B3;
defparam prom_inst_0.INIT_RAM_0D = 256'hECECEBEBEAE9E9E8E7E7E6E5E4E4E3E2E1E1E0DFDEDEDDDCDBDAD9D8D7D6D5D4;
defparam prom_inst_0.INIT_RAM_0E = 256'hFBFBFBFAFAF9F9F9F8F8F8F7F7F6F6F5F5F5F4F4F3F3F2F2F1F1F0EFEFEEEEED;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEFEFEFEFEFDFDFDFDFCFCFCFB;
defparam prom_inst_0.INIT_RAM_10 = 256'hFBFBFCFCFCFCFDFDFDFDFEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hECEDEDEEEFEFF0F0F1F1F2F2F3F3F4F4F5F5F6F6F7F7F7F8F8F9F9F9FAFAFAFB;
defparam prom_inst_0.INIT_RAM_12 = 256'hD4D5D5D6D7D8D9DADBDBDCDDDEDFE0E0E1E2E3E3E4E5E6E6E7E8E8E9EAEAEBEC;
defparam prom_inst_0.INIT_RAM_13 = 256'hB2B3B4B5B6B8B9BABBBCBDBEBFC1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3;
defparam prom_inst_0.INIT_RAM_14 = 256'h87888A8B8C8E8F919294959698999B9C9D9FA0A1A3A4A5A6A8A9AAACADAEAFB0;
defparam prom_inst_0.INIT_RAM_15 = 256'h535556585A5B5D5F6162646667696B6C6E6F7173747677797A7C7E7F81828485;
defparam prom_inst_0.INIT_RAM_16 = 256'h17191B1D1F21232527292A2C2E30323436383A3B3D3F41434546484A4C4E4F51;
defparam prom_inst_0.INIT_RAM_17 = 256'hD3D5D8DADCDEE0E3E5E7E9EBEDF0F2F4F6F8FAFCFE00030507090B0D0F111315;
defparam prom_inst_0.INIT_RAM_18 = 256'h898B8E909295979A9C9EA1A3A5A8AAACAFB1B3B6B8BABDBFC1C4C6C8CACDCFD1;
defparam prom_inst_0.INIT_RAM_19 = 256'h383A3D404245474A4D4F525457595C5E616466696B6E707375777A7C7F818486;
defparam prom_inst_0.INIT_RAM_1A = 256'hE2E4E7EAEDEFF2F5F8FAFD000205080B0D101315181B1D202325282B2D303335;
defparam prom_inst_0.INIT_RAM_1B = 256'h878A8C8F9295989B9EA1A3A6A9ACAFB2B5B7BABDC0C3C6C8CBCED1D4D6D9DCDF;
defparam prom_inst_0.INIT_RAM_1C = 256'h282B2E3134373A3D404346494C4F5255585B5E616366696C6F7275787B7E8184;
defparam prom_inst_0.INIT_RAM_1D = 256'hC6C9CCD0D3D6D9DCDFE2E5E8EBEEF1F4F7FAFE0104070A0D101316191C1F2225;
defparam prom_inst_0.INIT_RAM_1E = 256'h6366696C6F7276797C7F8285888B8F9295989B9EA1A4A7ABAEB1B4B7BABDC0C3;
defparam prom_inst_0.INIT_RAM_1F = 256'hFE0205080B0E1114181B1E2124272A2E3134373A3D4044474A4D505356595D60;
defparam prom_inst_0.INIT_RAM_20 = 256'h9A9DA0A3A7AAADB0B3B6B9BCC0C3C6C9CCCFD2D6D9DCDFE2E5E8ECEFF2F5F8FB;
defparam prom_inst_0.INIT_RAM_21 = 256'h373A3D404346494C4F5255595C5F6265686B6E7175787B7E8184878A8E919497;
defparam prom_inst_0.INIT_RAM_22 = 256'hD5D8DBDEE1E4E7EAEDF0F3F6F9FCFF0206090C0F1215181B1E2124272A2D3034;
defparam prom_inst_0.INIT_RAM_23 = 256'h76797C7F8285888B8E9194979A9D9FA2A5A8ABAEB1B4B7BABDC0C3C6C9CCCFD2;
defparam prom_inst_0.INIT_RAM_24 = 256'h1C1E2124272A2C2F3235383A3D404346494B4E5154575A5D5F6265686B6E7174;
defparam prom_inst_0.INIT_RAM_25 = 256'hC6C8CBCDD0D3D5D8DBDDE0E3E5E8EBEDF0F3F5F8FBFE000306080B0E11131619;
defparam prom_inst_0.INIT_RAM_26 = 256'h75777A7C7F818486898B8D909295979A9C9FA2A4A7A9ACAEB1B3B6B9BBBEC0C3;
defparam prom_inst_0.INIT_RAM_27 = 256'h2B2D2F313336383A3C3F414346484A4D4F515456585B5D5F626466696B6E7072;
defparam prom_inst_0.INIT_RAM_28 = 256'hE7E9EBEDEFF1F3F5F7F9FBFD00020406080A0C0E10131517191B1D2022242628;
defparam prom_inst_0.INIT_RAM_29 = 256'hABADAFB1B2B4B6B8BABBBDBFC1C3C5C6C8CACCCED0D2D4D6D7D9DBDDDFE1E3E5;
defparam prom_inst_0.INIT_RAM_2A = 256'h78797B7C7E7F8182848687898A8C8D8F9192949597999A9C9E9FA1A3A5A6A8AA;
defparam prom_inst_0.INIT_RAM_2B = 256'h4D4E50515253545657585A5B5C5D5F606163646567686A6B6C6E6F7172747576;
defparam prom_inst_0.INIT_RAM_2C = 256'h2B2C2D2E2F303132333435363738393A3B3C3D3E3F41424344454647484A4B4C;
defparam prom_inst_0.INIT_RAM_2D = 256'h131414151616171818191A1A1B1C1D1D1E1F2020212223242525262728292A2B;
defparam prom_inst_0.INIT_RAM_2E = 256'h05050506060607070708080909090A0A0B0B0C0C0D0D0E0E0F0F101011111213;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000000000000000000000010101010101010102020202020303030304040404;
defparam prom_inst_0.INIT_RAM_30 = 256'h0505050404040303030302020202020201010101010101000000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h14141312121111100F0F0E0E0D0D0C0C0B0B0B0A0A0909080808070707060605;
defparam prom_inst_0.INIT_RAM_32 = 256'h2D2C2B2A2928272726252423222221201F1F1E1D1C1C1B1A1919181717161515;
defparam prom_inst_0.INIT_RAM_33 = 256'h4F4E4D4B4A4948474644434241403F3E3D3C3B3A393736353433333231302F2E;
defparam prom_inst_0.INIT_RAM_34 = 256'h7A797776747371706F6D6C6A696866656362615F5E5D5B5A5958565554535150;
defparam prom_inst_0.INIT_RAM_35 = 256'hAEACABA9A7A5A4A2A09F9D9B9A9896959391908E8D8B898886858382807F7D7C;
defparam prom_inst_0.INIT_RAM_36 = 256'hEAE8E6E4E2E0DEDCDAD8D7D5D3D1CFCDCBC9C7C6C4C2C0BEBCBBB9B7B5B3B2B0;
defparam prom_inst_0.INIT_RAM_37 = 256'h2E2C29272523211E1C1A181614110F0D0B0907050301FFFCFAF8F6F4F2F0EEEC;
defparam prom_inst_0.INIT_RAM_38 = 256'h797674716F6C6A686563615E5C59575552504E4B49474442403E3B3937353230;
defparam prom_inst_0.INIT_RAM_39 = 256'hC9C7C4C2BFBCBAB7B5B2B0ADAAA8A5A3A09E9B999694918F8C8A878582807D7B;
defparam prom_inst_0.INIT_RAM_3A = 256'h201D1A1815120F0D0A070402FFFCF9F7F4F1EFECE9E7E4E1DFDCD9D7D4D1CFCC;
defparam prom_inst_0.INIT_RAM_3B = 256'h7B7875726F6C696764615E5B585553504D4A4744413F3C393633312E2B282523;
defparam prom_inst_0.INIT_RAM_3C = 256'hDAD7D4D1CECBC8C5C2BFBCB9B6B3B0ADAAA7A4A19E9B9895928F8C898784817E;
defparam prom_inst_0.INIT_RAM_3D = 256'h3B3835322F2C292623201C191613100D0A070401FEFBF8F5F2EFECE9E6E3E0DD;
defparam prom_inst_0.INIT_RAM_3E = 256'h9F9C9895928F8C8986837F7C797673706D6A6763605D5A5754514E4B4844413E;
defparam prom_inst_0.INIT_RAM_3F = 256'h0300FDFAF7F3F0EDEAE7E4E1DDDAD7D4D1CECBC7C4C1BEBBB8B5B1AEABA8A5A2;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[28:0],dout[10:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[10:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h4444444444444444444444444444444444444444444444444444444444444444;
defparam prom_inst_1.INIT_RAM_01 = 256'h5555555555555555555555555555555555555555555555444444444444444444;
defparam prom_inst_1.INIT_RAM_02 = 256'h6666666666666666666666555555555555555555555555555555555555555555;
defparam prom_inst_1.INIT_RAM_03 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam prom_inst_1.INIT_RAM_04 = 256'h7777777777777777777777777777777777777777777766666666666666666666;
defparam prom_inst_1.INIT_RAM_05 = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_06 = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_07 = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_08 = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_09 = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_0A = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_0B = 256'h6666666666666666666667777777777777777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_0C = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam prom_inst_1.INIT_RAM_0D = 256'h5555555555555555555555555555555555555555555666666666666666666666;
defparam prom_inst_1.INIT_RAM_0E = 256'h4444444444444444444555555555555555555555555555555555555555555555;
defparam prom_inst_1.INIT_RAM_0F = 256'h3444444444444444444444444444444444444444444444444444444444444444;
defparam prom_inst_1.INIT_RAM_10 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam prom_inst_1.INIT_RAM_11 = 256'h2222222222222222222222222222222222222222222222233333333333333333;
defparam prom_inst_1.INIT_RAM_12 = 256'h1111111111111111111111222222222222222222222222222222222222222222;
defparam prom_inst_1.INIT_RAM_13 = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam prom_inst_1.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000011111111111111111111;
defparam prom_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h1111111111111111111111000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam prom_inst_1.INIT_RAM_1D = 256'h2222222222222222222222222222222222222222222211111111111111111111;
defparam prom_inst_1.INIT_RAM_1E = 256'h3333333333333333333322222222222222222222222222222222222222222222;
defparam prom_inst_1.INIT_RAM_1F = 256'h4433333333333333333333333333333333333333333333333333333333333333;

endmodule //Gowin_pROM
