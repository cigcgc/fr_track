parameter INTEGER_WIDTH = 16;
