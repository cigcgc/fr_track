parameter NUM_CHN=1;
parameter DATA_WIDTH=16;
parameter PARAM_FRACTION_WIDTH=8;
