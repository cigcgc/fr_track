`define MODULE_NAME Fixed_to_Float_Top
`define NO_CE
`define Custom
