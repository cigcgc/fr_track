`define MODULE_NAME PID_Controller_3p3z_Top
